module moduleName (
    input a
);
    
endmodule